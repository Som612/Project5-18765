   `celldefine
module scanff(CK, SD, SI, SE, Q);
    input CK, SD, SI, SE, Q;
    output Q;

    wire a;
    sff(Q, CK, a);
    u_mux2 (a, SD, SI, SE);

endmodule
`endcelldefine

module s9234_scan(Din, scan_in, SE, Clk, scan_out, g89,g94,g98,g102,g107,g301,g306,g310,g314,g319,g557,g558,g559,g560,g561,
  g562,g563,g564,g705,g639,g567,g45,g42,g39,g702,g32,g38,g46,g36,g47,g40,g37,
  g41,g22,g44,g23,g678,g332,g123,g207,g695,g461,g18, g292,g331,g689,g24,g465,g84,g291,g676,g622,g117,g278,g128,
  g598,g554,g496,g179,g48,g590,g551,g682,g11,g606,g188,g646,g327,g361,g289,g398,g684,g619,g208,g248,g390,g625,
  g681,g437,g276,g3,g323,g224,g685,g43,g157,g282,g697,g206,g449,g118,g528,g284,g426,g634,g669,g520,g281,g175,g15,
  g631,g69,g693,g337,g457,g486,g471,g328,g285,g418,g402,g297,g212,g410,g430,g33,g662,g453,g269,g574,g441,g664,
  g349,g211,g586,g571,g29,g326,g698,g654,g293,g690,g445,g374,g6,g687,g357,g386,g504,g665,g166,g541,g74,g338,g696,
  g516,g536,g683,g353,g545,g254,g341,g290,g2,g287,g336,g345,g628,g679,g28,g688,g283,g613,g10,g14,g680,g143,g672,
  g667,g366,g279,g492,g170,g686,g288,g638,g602,g642,g280,g663,g610,g148,g209,g675,g478,g122,g54,g594,g286,g616,g79,
  g218,g242,g578,g184,g119,g668,g139,g422,g210,g394,g230,g25,g204,g658,g650,g378,g508,g548,g370,g406,g236,g500,g205,
  g197,g666,g114,g524,g260,g111,g131,g7,g19,g677,g582,g485,g699,g193,g135,g382,g414,g434,g266,g49,g152,g692,g277,
  g127,g161,g512,g532,g64,g694,g691,g1,g59,g2584,g3222,g3600,g4307,g4321,g4422,g4809,g5137,g5468,g5469,g5692,g6282,
  g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,g6374,g6728,g1290,g4121,g4108,g4106,g4103,g1293,g4099,g4102,g4109,
  g4100,g4112,g4105,g4101,g4110,g4104,g4107,g4098,g4130,g6823,g6940,g6102,g4147,g4841,g6725,g3232,g4119,g4141,g6726,
  g6507,g6590,g3231,g5330,g5147,g4839,g6105,g5138,g4122,g6827,g6745,g6405,g6729,g6595,g6826,g4134,g6599,g4857,g6406,
  g5148,g4117,g6582,g3229,g5700,g4136,g4858,g5876,g3239,g5698,g5328,g4133,g4847,g5877,g6597,g4120,g3235,g4137,g6407,
  g5470,g6841,g4149,g6101,g4844,g4113,g6504,g3224,g4855,g4424,g5582,g6502,g6107,g5472,g6602,g5581,g6587,g4145,g2585,
  g4842,g2586,g1291,g4118,g3225,g4853,g4849,g6512,g3233,g4851,g4856,g6854,g1831,g4843,g6510,g6591,g4846,g1288,g5478,
  g6840,g6594,g5580,g6853,g4840,g4150,g5490,g6511,g4142,g4845,g5694,g6722,g4139,g5480,g5697,g6498,g4126,g5471,g6505,
  g6588,g5475,g4148,g6501,g6506,g4135,g5476,g3230,g6721,g3227,g6925,g5477,g5489,g4131,g6727,g4140,g6842,g4423,g6723,
  g6724,g4132,g6401,g5491,g4127,g6278,g6106,g6744,g6404,g4138,g3228,g1289,g4123,g4658,g5878,g4125,g4124,g5874,g6103,
  g1294,g1292,g4115,g6584,g6596,g3226,g2587,g4657,g6589,g3234,g3238,g6592,g5473,g4114,g6800,g5141,g4854,g6839,g5695,
  g6499,g6825,g5693,g4850,g3237,g6497,g6100,g6509,g4128,g4116,g6503,g3241,g489);

  input Din, scan_in, SE, Clk, g89,g94,g98,g102,g107,g301,g306,g310,g314,g319,g557,g558,g559,g560,g561,
  g562,g563,g564,g705,g639,g567,g45,g42,g39,g702,g32,g38,g46,g36,g47,g40,g37,
  g41,g22,g44,g23,g678,g332,g123,g207,g695,g461,g18, g292,g331,g689,g24,g465,g84,g291,g676,g622,g117,g278,g128,
  g598,g554,g496,g179,g48,g590,g551,g682,g11,g606,g188,g646,g327,g361,g289,g398,g684,g619,g208,g248,g390,g625,
  g681,g437,g276,g3,g323,g224,g685,g43,g157,g282,g697,g206,g449,g118,g528,g284,g426,g634,g669,g520,g281,g175,
  g15,g631,g69,g693,g337,g457,g486,g471,g328,g285,g418,g402,g297,g212,g410,g430,g33,g662,g453,g269,g574,g441,g664,
  g349,g211,g586,g571,g29,g326,g698,g654,g293,g690,g445,g374,g6,g687,g357,g386,g504,g665,g166,g541,g74,g338,g696,
  g516,g536,g683,g353,g545,g254,g341,g290,g2,g287,g336,g345,g628,g679,g28,g688,g283,g613,g10,g14,g680,g143,g672,
  g667,g366,g279,g492,g170,g686,g288,g638,g602,g642,g280,g663,g610,g148,g209,g675,g478,g122,g54,g594,g286,g616,g79,
  g218,g242,g578,g184,g119,g668,g139,g422,g210,g394,g230,g25,g204,g658,g650,g378,g508,g548,g370,g406,g236,g500,g205,
  g197,g666,g114,g524,g260,g111,g131,g7,g19,g677,g582,g485,g699,g193,g135,g382,g414,g434,g266,g49,g152,g692,g277,
  g127,g161,g512,g532,g64,g694,g691,g1,g59,g489;

  output scan_out,g2584,g3222,g3600,g4307,g4321,g4422,g4809,g5137,g5468,g5469,g5692,g6282,g6284,g6360,g6362,g6364,g6366,
  g6368,g6370,g6372,g6374,g6728,g1290,g4121,g4108,g4106,g4103,g1293,g4099,g4102,g4109,g4100,g4112,g4105,g4101,g4110,
  g4104,g4107,g4098,g4130,g6823,g6940,g6102,g4147,g4841,g6725,g3232,g4119,g4141,g6726,g6507,g6590,g3231,g5330,g5147,
  g4839,g6105,g5138,g4122,g6827,g6745,g6405,g6729,g6595,g6826,g4134,g6599,g4857,g6406,g5148,g4117,g6582,g3229,g5700,  
  g4136,g4858,g5876,g3239,g5698,g5328,g4133,g4847,g5877,g6597,g4120,g3235,g4137,g6407,g5470,g6841,g4149,g6101,g4844,  
  g4113,g6504,g3224,g4855,g4424,g5582,g6502,g6107,g5472,g6602,g5581,g6587,g4145,g2585,g4842,g2586,g1291,g4118,g3225,
  g4853,g4849,g6512,g3233,g4851,g4856,g6854,g1831,g4843,g6510,g6591,g4846,g1288,g5478,g6840,g6594,g5580,g6853,g4840,
  g4150,g5490,g6511,g4142,g4845,g5694,g6722,g4139,g5480,g5697,g6498,g4126,g5471,g6505,g6588,g5475,g4148,g6501,g6506,
  g4135,g5476,g3230,g6721,g3227,g6925,g5477,g5489,g4131,g6727,g4140,g6842,g4423,g6723,g6724,  g4132,g6401,g5491,g4127,
  g6278,g6106,g6744,g6404,g4138,g3228,g1289,g4123,g4658,g5878,g4125,g4124,g5874,g6103,g1294,g1292,g4115,g6584,g6596,
  g3226,g2587,g4657,g6589,g3234,g3238,g6592,g5473,g4114,g6800,g5141,g4854,g6839,g5695,  g6499,g6825,g5693,g4850,g3237,
  g6497,g6100,g6509,g4128,g4116,g6503,g3241;

  wire g678, g332, g6940,g6102,g4147,g4841,g6725,g3232,g4119,g4141,g6726,g6507,g6590,g3231,g5330,g5147,g4839,g6105,g5138,
  g4122,g6827,g6745,g6405,g6729,g6595,g6826,g4134,g6599,g4857,g6406,g5148,g4117,g6582,g3229,g5700,g4136,g4858,g5876,g3239,
  g5698,g5328,g4133,g4847,g5877,g6597,g4120,g3235,g4137,g6407,g5470,g6841,g4149,g6101,g4844,g4113,g6504,g3224,g4855,g4424,
  g5582,g6502,g6107,g5472,g6602,g5581,g6587,g4145,g2585,g4842,g2586,g1291,g4118,g3225,g4853,g4849,g6512,g3233,g4851,g4856,
  g6854,g1831,g4843,g6510,g6591,g4846,g1288,g5478,g6840,g6594,g5580,g6853,g4840,g4150,g5490,g6511,g4142,g4845,g5694,g6722,
  g4139,g5480,g5697,g6498,g4126,g5471,g6505,g6588,g5475,g4148,g6501,g6506,g4135,g5479,g6824,g3240,g5476,g3230,g6721,g3227,
  g6925,g5477,g5489,g4131,g6727,g4140,g6842,g4423,g6723,g6724,g4132,g6401,g5491,g4127,g6278,g6106,g6744,g6404,g4138,g3228,
  g1289,g4123,g4658,g5878,g4125,g4124,g5874,g6103,g1294,g1292,g4115,g6584,g6596,g3226,g2587,g4657,g6589,g3234,g3238,g6592,
  g5473,g4114,g6800,g5241,g4584,g6839,g5699,g3236,g6601,g5875,g4425,g5329,g5695,g6499,g6825,g5693,g4850,g3237,g6497,g6100,
  g6509,g4128,g4116,g6503,g3241,g6277,g5139,g6598,g6600,g4129,g6593,g6801,g4426,g5474,g5140,g5696,g4852,g4848,g4659,g6583,
  g6402,g4144,g6104,g6941,g6403,g6500,g6508,g6586,g4146,g4143,g6720,g6585;


  sff SFF_0(CK,g4130,scan_in,SE,g678);
  sff SFF_1(CK,g6823,g678,SE,g332);
  sff SFF_2(CK,g123,g332,SE,g6940);
  sff SFF_3(CK,g207,g6940,SE,g6102);
  sff SFF_4(CK,g695,g6102,SE,g4147);
  sff SFF_5(CK,g461,g4147,SE,g4841);
  sff SFF_6(CK,g18,g4841,SE,g6725);
  sff SFF_7(CK,g292,g6725,SE,g3232);
  sff SFF_8(CK,g331,g3232,SE,g4119);
  sff SFF_9(CK,g689,g4119,SE,g4141);
  sff SFF_10(CK,g24,g4141,SE,g6726);
  sff SFF_11(CK,g465,g6726,SE,g6507);
  sff SFF_12(CK,g84,g6507,SE,g6590);
  sff SFF_13(CK,g291,g6590,SE,g3231);
  sff SFF_14(CK,g676,g3231,SE,g5330);
  sff SFF_15(CK,g622,g5330,SE,g5147);
  sff SFF_16(CK,g117,g5147,SE,g4839);
  sff SFF_17(CK,g278,g839,SE,g6105);
  sff SFF_18(CK,g128,g6105,SE,g5138);
  sff SFF_19(CK,g598,g5138,SE,g4122);
  sff SFF_20(CK,g554,g4122,SE,g6827);
  sff SFF_21(CK,g496,g6827,SE,g6745);
  sff SFF_22(CK,g179,g6745,SE,g6405);
  sff SFF_23(CK,g48,g6405,SE,g6729);
  sff SFF_24(CK,g590,g6729,SE,g6595);
  sff SFF_25(CK,g551,g6595,SE,g6826);
  sff SFF_26(CK,g682,g6826,SE,g4134);
  sff SFF_27(CK,g11,g4134,SE,g6599);
  sff SFF_28(CK,g606,g6599,SE,g4857);
  sff SFF_29(CK,g188,g4857,SE,g6406);
  sff SFF_30(CK,g646,g6406,SE,g5148);
  sff SFF_31(CK,g327,g5148,SE,g4117);
  sff SFF_32(CK,g361,g4117,SE,g6582);
  sff SFF_33(CK,g289,g6582,SE,g3229);
  sff SFF_34(CK,g398,g3229,SE,g5700);
  sff SFF_35(CK,g684,g5700,SE,g4136);
  sff SFF_36(CK,g619,g4136,SE,g4858);
  sff SFF_37(CK,g208,g4858,SE,g5876);
  sff SFF_38(CK,g248,g5876,SE,g3239);
  sff SFF_39(CK,g390,g3239,SE,g5698);
  sff SFF_40(CK,g625,g5698,SE,g5328);
  sff SFF_41(CK,g681,g5328,SE,g4133);
  sff SFF_42(CK,g437,g4133,SE,g4847);
  sff SFF_43(CK,g276,g4847,SE,g5877);
  sff SFF_44(CK,g3,g5877,SE,g6597);
  sff SFF_45(CK,g323,g6597,SE,g4120);
  sff SFF_46(CK,g224,g4120,SE,g3235);
  sff SFF_47(CK,g685,g3235,SE,g4137);
  sff SFF_48(CK,g43,g4137,SE,g6407);
  sff SFF_49(CK,g157,g6407,SE,g5470);
  sff SFF_50(CK,g282,g5470,SE,g6841);
  sff SFF_51(CK,g697,g6841,SE,g4149);
  sff SFF_52(CK,g206,g4149,SE,g6101);
  sff SFF_53(CK,g449,g6101,SE,g4844);
  sff SFF_54(CK,g118,g4844,SE,g4113);
  sff SFF_55(CK,g528,g4113,SE,g6504);
  sff SFF_56(CK,g284,g6504,SE,g3224);
  sff SFF_57(CK,g426,g3224,SE,g4855);
  sff SFF_58(CK,g634,g4855,SE,g4424);
  sff SFF_59(CK,g669,g4424,SE,g5582);
  sff SFF_60(CK,g520,g5582,SE,g6502);
  sff SFF_61(CK,g281,g6502,SE,g6107);
  sff SFF_62(CK,g175,g6107,SE,g5472);
  sff SFF_63(CK,g15,g5472,SE,g6602);
  sff SFF_64(CK,g631,g6602,SE,g5581);
  sff SFF_65(CK,g69,g5581,SE,g6587);
  sff SFF_66(CK,g693,g6587,SE,g4145);
  sff SFF_67(CK,g337,g4145,SE,g2585);
  sff SFF_68(CK,g457,g2585,SE,g4842);
  sff SFF_69(CK,g486,g4842,SE,g2586);
  sff SFF_70(CK,g471,g2586,SE,g1291);
  sff SFF_71(CK,g328,g1291,SE,g4118);
  sff SFF_72(CK,g285,g4118,SE,g3225);
  sff SFF_73(CK,g418,g3225,SE,g4853);
  sff SFF_74(CK,g402,g4853,SE,g4849);
  sff SFF_75(CK,g297,g4849,SE,g6512);
  sff SFF_76(CK,g212,g6512,SE,g3233);
  sff SFF_77(CK,g410,g3233,SE,g4851);
  sff SFF_78(CK,g430,g4851,SE,g4856);
  sff SFF_79(CK,g33,g4856,SE,g6854);
  sff SFF_80(CK,g662,g6854,SE,g1831);
  sff SFF_81(CK,g453,g1831,SE,g4843);
  sff SFF_82(CK,g269,g4843,SE,g6510);
  sff SFF_83(CK,g574,g6510,SE,g6591);
  sff SFF_84(CK,g441,g6591,SE,g4846);
  sff SFF_85(CK,g664,g4846,SE,g1288);
  sff SFF_86(CK,g349,g1288,SE,g5478);
  sff SFF_87(CK,g211,g5478,SE,g6840);
  sff SFF_88(CK,g586,g6840,SE,g6594);
  sff SFF_89(CK,g571,g6594,SE,g5580);
  sff SFF_90(CK,g29,g5580,SE,g6853);
  sff SFF_91(CK,g326,g6853,SE,g4840);
  sff SFF_92(CK,g698,g4840,SE,g4150);
  sff SFF_93(CK,g654,g4150,SE,g5490);
  sff SFF_94(CK,g293,g5490,SE,g6511);
  sff SFF_95(CK,g690,g6511,SE,g4142);
  sff SFF_96(CK,g445,g4142,SE,g4845);
  sff SFF_97(CK,g374,g4845,SE,g5694);
  sff SFF_98(CK,g6,g5694,SE,g6722);
  sff SFF_99(CK,g687,g6722,SE,g4139);
  sff SFF_100(CK,g357,g4139,SE,g5480);
  sff SFF_101(CK,g386,g5480,SE,g5697);
  sff SFF_102(CK,g504,g5697,SE,g6498);
  sff SFF_103(CK,g665,g6498,SE,g4126);
  sff SFF_104(CK,g166,g4126,SE,g5471);
  sff SFF_105(CK,g541,g5471,SE,g6505);
  sff SFF_106(CK,g74,g6505,SE,g6588);
  sff SFF_107(CK,g338,g6588,SE,g5475);
  sff SFF_108(CK,g696,g5475,SE,g4148);
  sff SFF_109(CK,g516,g4148,SE,g6501);
  sff SFF_110(CK,g536,g6501,SE,g6506);
  sff SFF_111(CK,g683,g6506,SE,g4135);
  sff SFF_112(CK,g353,g4135,SE,g5479);
  sff SFF_113(CK,g545,g5479,SE,g6824);
  sff SFF_114(CK,g254,g6824,SE,g3240);
  sff SFF_115(CK,g341,g3240,SE,g5476);
  sff SFF_116(CK,g290,g5476,SE,g3230);
  sff SFF_117(CK,g2,g3230,SE,g6721);
  sff SFF_118(CK,g287,g6721,SE,g3227);
  sff SFF_119(CK,g336,g3227,SE,g6925);
  sff SFF_120(CK,g345,g6925,SE,g5477);
  sff SFF_121(CK,g628,g5477,SE,g5489);
  sff SFF_122(CK,g679,g5489,SE,g4131);
  sff SFF_123(CK,g28,g4131,SE,g6727);
  sff SFF_124(CK,g688,g6727,SE,g4140);
  sff SFF_125(CK,g283,g4140,SE,g6842);
  sff SFF_126(CK,g613,g6842,SE,g4423);
  sff SFF_127(CK,g10,g4423,SE,g6723);
  sff SFF_128(CK,g14,g6723,SE,g6724);
  sff SFF_129(CK,g680,g6724,SE,g4132);
  sff SFF_130(CK,g143,g4132,SE,g6401);
  sff SFF_131(CK,g672,g6401,SE,g5491);
  sff SFF_132(CK,g667,g5491,SE,g4127);
  sff SFF_133(CK,g366,g4127,SE,g6278);
  sff SFF_134(CK,g279,g6278,SE,g6106);
  sff SFF_135(CK,g492,g6106,SE,g6744);
  sff SFF_136(CK,g170,g6744,SE,g6404);
  sff SFF_137(CK,g686,g6404,SE,g4138);
  sff SFF_138(CK,g288,g4138,SE,g3228);
  sff SFF_139(CK,g638,g3228,SE,g1289);
  sff SFF_140(CK,g602,g1289,SE,g4123);
  sff SFF_141(CK,g642,g4123,SE,g4658);
  sff SFF_142(CK,g280,g4658,SE,g5878);
  sff SFF_143(CK,g663,g5878,SE,g4125);
  sff SFF_144(CK,g610,g4125,SE,g4124);
  sff SFF_145(CK,g148,g4124,SE,g5874);
  sff SFF_146(CK,g209,g5874,SE,g6103);
  sff SFF_147(CK,g675,g6103,SE,g1294);
  sff SFF_148(CK,g478,g1294,SE,g1292);
  sff SFF_149(CK,g122,g1292,SE,g4115);
  sff SFF_150(CK,g54,g4115,SE,g6584);
  sff SFF_151(CK,g594,g6584,SE,g6596);
  sff SFF_152(CK,g286,g6596,SE,g3226);
  sff SFF_153(CK,g489,g3226,SE,g2587);
  sff SFF_154(CK,g616,g2587,SE,g4657);
  sff SFF_155(CK,g79,g4657,SE,g6589);
  sff SFF_156(CK,g218,g6589,SE,g3234);
  sff SFF_157(CK,g242,g3234,SE,g3238);
  sff SFF_158(CK,g578,g3238,SE,g6592);
  sff SFF_159(CK,g184,g6592,SE,g5473);
  sff SFF_160(CK,g119,g5473,SE,g4114);
  sff SFF_161(CK,g668,g4114,SE,g6800);
  sff SFF_162(CK,g139,g6800,SE,g5141);
  sff SFF_163(CK,g422,g5141,SE,g4854);
  sff SFF_164(CK,g210,g4854,SE,g6839);
  sff SFF_165(CK,g394,g6839,SE,g5699);
  sff SFF_166(CK,g230,g5699,SE,g3236);
  sff SFF_167(CK,g25,g3236,SE,g6601);
  sff SFF_168(CK,g204,g6601,SE,g5875);
  sff SFF_169(CK,g658,g5875,SE,g4425);
  sff SFF_170(CK,g650,g4425,SE,g5329);
  sff SFF_171(CK,g378,g5329,SE,g5695);
  sff SFF_172(CK,g508,g5695,SE,g6499);
  sff SFF_173(CK,g548,g6499,SE,g6825);
  sff SFF_174(CK,g370,g6825,SE,g5693);
  sff SFF_175(CK,g406,g6593,SE,g4850);
  sff SFF_176(CK,g236,g4850,SE,g3237);
  sff SFF_177(CK,g500,g3237,SE,g6497);
  sff SFF_178(CK,g205,g6497,SE,g6100);
  sff SFF_179(CK,g197,g6100,SE,g6509);
  sff SFF_180(CK,g666,g6509,SE,g4128);
  sff SFF_181(CK,g114,g4128,SE,g4116);
  sff SFF_182(CK,g524,g4116,SE,g6503);
  sff SFF_183(CK,g260,g6503,SE,g3241);
  sff SFF_184(CK,g111,g3241,SE,g6277);
  sff SFF_185(CK,g131,g6277,SE,g5139);
  sff SFF_186(CK,g7,g5139,SE,g6598);
  sff SFF_187(CK,g19,g6598,SE,g6600);
  sff SFF_188(CK,g677,g6600,SE,g4129);
  sff SFF_189(CK,g582,g4129,SE,g6593);
  sff SFF_190(CK,g485,g6593,SE,g6801);
  sff SFF_191(CK,g699,g6801,SE,g4426);
  sff SFF_192(CK,g193,g4426,SE,g5474);
  sff SFF_193(CK,g135,g5474,SE,g5140);
  sff SFF_194(CK,g382,g5410,SE,g5696);
  sff SFF_195(CK,g414,g5696,SE,g4852);
  sff SFF_196(CK,g434,g4852,SE,g4848);
  sff SFF_197(CK,g266,g4848,SE,g4659);
  sff SFF_198(CK,g49,g4659,SE,g6583);
  sff SFF_199(CK,g152,g6583,SE,g6402);
  sff SFF_200(CK,g692,g6402,SE,g4144);
  sff SFF_201(CK,g277,g4144,SE,g6104);
  sff SFF_202(CK,g127,g6104,SE,g6941);
  sff SFF_203(CK,g161,g6941,SE,g6403);
  sff SFF_204(CK,g512,g6403,SE,g6500);
  sff SFF_205(CK,g532,g6500,SE,g6508);
  sff SFF_206(CK,g64,g6508,SE,g6586);
  sff SFF_207(CK,g694,g6586,SE,g4146);
  sff SFF_208(CK,g691,g4146,SE,g4143);
  sff SFF_209(CK,g1,g4143,SE,g6720);
  sff SFF_210(CK,g59,g6720,SE,scan_out);
  
endmodule






 

