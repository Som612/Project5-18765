//Large wrapper for Project 5
//Extra inputs for TAP: 4
//Extra inputs for instructions: 4
//Extra outputs for testing: 0,?

module DFT_full(data_in,data_out,clk,reset);

//Ports
input clk,reset;	//Clock input
input [44:0] data_in;//Inputs for the tap controller and circuit
output [38:0] data_out;//Response

//Wires

//Code Starts Here

endmodule//End of DFT Module

//4 to 1 MUX